module ForwardUnit(
    input Ex_Mem_RegWrite
)